cdl_package CYGPKG_DEVS_ETH_ARM_GALOIS {
    display       "Marvell ethernet driver for Galois SoC"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_ARM_ARM9_GALOIS

    include_dir   .
    include_files ; # none _exported_ whatsoever

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0

    description   "Ethernet driver for Marvell Galois SoC."
    compile       -library=libextras.a ethernet.c

    cdl_option CYGNUM_DEVS_ETH_ARM_GALOIS_CPUINDEX {
        display "Ethernet runs on CPU#0 or CPU#1"
        flavor  data
	legal_values 0 to 1
        default_value 0
        description "Ethernet runs on CPU#0 or CPU#1"
    }

    cdl_option CYGNUM_DEVS_ETH_ARM_GALOIS_TXQLEN {
        display       "Length of tx queue"
        flavor        data
        legal_values  2 to 128
        default_value 64
        description   "Length of tx queue"
    }

    cdl_option CYGNUM_DEVS_ETH_ARM_GALOIS_RXQLEN {
        display       "Length of rx queue"
        flavor        data
        legal_values  2 to 128
        default_value 64
        description   "Length of rx queue"
    }

    cdl_component CYGSEM_DEVS_ETH_ARM_GALOIS_2BSTUFF {
        display "2B stuff to rx packets"
        flavor  bool
        default_value 1
        description "2B stuff, see datasheet."
    }

    cdl_component CYGSEM_DEVS_ETH_ARM_GALOIS_10M {
        display "Fixed to 10Mb/s"
        flavor  bool
        default_value 1
        description "Fixed to 10Mb/s"
    }

    cdl_component CYGPKG_DEVS_ETH_ARM_GALOIS_OPTIONS {
        display "Galois ethernet driver build options"
        flavor  none
	    no_define

        cdl_option CYGPKG_DEVS_ETH_ARM_GALOIS_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Galois ethernet driver package. 
		        These flags are used in addition to the set of global 
		        flags."
        }
    }

}
