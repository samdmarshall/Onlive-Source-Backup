# ====================================================================
#
#      hal_coldfire_m5272c3.cdl
#
#      Freescale M5272C3 evaluation board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2006 eCosCentric Ltd.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):     Enrico Piria
## Contributors:  Wade Jensen
## Date:          2005-25-06
##
######DESCRIPTIONEND####
##========================================================================

cdl_package CYGPKG_HAL_COLDFIRE_M5272C3 {
    display         "Freescale M5272C3 evaluation board"
    parent          CYGPKG_HAL_COLDFIRE_MCF5272
    define_header   hal_coldfire_m5272c3.h
    include_dir     cyg/hal

    description   "The Freescale M5272C3 evaluation board platform HAL
                package should be used when targeting the actual hardware for
                the Freescale M5272C3 evaluation board platform."

    compile     plf_startup.c

    implements      CYGINT_HAL_DEBUG_GDB_STUBS
    implements      CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements      CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT


    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_coldfire.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_coldfire_mcf5272.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_coldfire_m5272c3.h>"
        puts $::cdl_system_header "#define HAL_PLATFORM_BOARD    \"Freescale M5272C3\""
        puts $::cdl_system_header "#define HAL_PLATFORM_EXTRA    \"\""
    }

    # The "-o file" is a workaround for CR100958 - without it the
    # output file would end up in the source directory under CygWin.
    # n.b. grep does not behave itself under win32
    make -priority 1 {
        <PREFIX>/include/cyg/hal/plf_offsets.inc : <PACKAGE>/src/plf_mk_defs.c
        $(CC) $(ACTUAL_CFLAGS) $(INCLUDE_PATH) -Wp,-MD,plf_offsets.tmp -o plf_mk_defs.tmp -S $<
        fgrep .equ plf_mk_defs.tmp | sed s/#// > $@
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 plf_offsets.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm plf_offsets.tmp plf_mk_defs.tmp
    }

    cdl_component CYG_HAL_STARTUP {
        display         "Startup type"
        flavor          data
        legal_values    {"RAM" "ROM" "ROMRAM"}
        default_value   {"RAM"}
        no_define
        define -file system.h CYG_HAL_STARTUP

        description "
           This option is used to control where the application program will
           run, either from RAM or ROM (flash) memory. ROM based applications
           must be self contained, while RAM applications will typically assume
           the existence of a debug environment, such as GDB stubs.
           ROMRAM bootstrap is similar to ROM bootstrap, but everything
           is copied to RAM before execution starts, thus improving performace,
           but at the cost of an increased RAM footprint."
    }
    
    cdl_option CYGHWR_HAL_ROM_LMA {
       display          "Load address for ROM image"
       active_if        { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "ROMRAM" }
       flavor           data
       legal_values     0xFFE00000 0xFFF00000
       default_value    0xFFF00000

       description    "This option lets you decide in which half of flash
                    memory to download the ROM image. As a safety measure,
                    the default is to use the upper half (starting at
                    0xFFF00000), thus preserving the ROM monitor shipped with
                    the board. This option is meaningful only when ROM or
                    ROMRAM startup is choosed."
    }
    
    cdl_option CYGHWR_HAL_SYSTEM_CLOCK_MHZ {
       display          "System clock speed in MHz"
       flavor           data
       legal_values     66 48
       default_value    66

       description    "This option identifies the system clock that the
                    processor uses. This value is used to set clock dividers
                    for some devices."
    }

    cdl_option CYGHWR_EXT_SRAM_INSTALLED {
       display          "External 512Kb SRAM module"
       flavor           bool
       default_value    0

       description    "If this option is enabled, chip-select module 2 is
           configured to access the optional external 512Kb SRAM module."
    }

    cdl_option CYGHWR_INSTALLED_SDRAM_SIZE {
       display          "Megabytes of SDRAM installed"
       flavor           data
       legal_values     16 4
       default_value    16

       description    "This option selects the size of the SDRAM installed.
            Note that the linker scripts have been written for a board with
            16 Mb of RAM. If you modify this option, you will have to change
            them by hand."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
       display          "Number of communication channels on the board"
       flavor           data
       calculated       2
       description      "
            Port 0 is the terminal serial port; port 1 is the auxiliary
            serial port."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
       display          "Debug serial port"
       active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
       flavor data
       legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
       default_value    0
       description      "
           This option chooses which port will be used to connect to a host
           via the GDB remote protocol."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "Debug serial port baud rate"
        active_if     CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 19200
        description   "
            This option controls the baud rate used for the GDB connection."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           This option chooses which port will be used for diagnostic output."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
       display          "Diagnostic serial port baud rate"
       active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
       flavor           data
       legal_values     9600 19200 38400 57600 115200
       default_value    19200

       description    "This option selects the baud rate used for the
                    diagnostic port. Note: this should match the value chosen
                    for the GDB port if the diagnostic and GDB port are the
                    same."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none

        description   "Set the periodic timer on the MCF5272 to 10 ms or
                    10000000 ns."

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value 4125
            description   "
                The default value is calculated as: 
                10 ms / ((1 / (66 MHz)) * 16 * 10)."
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE

        description   "Global build options including control over compiler
                    flags, linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "m68k-elf" }

            description       "This option specifies the command prefix used
                            when invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-m5206e -malign-int -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -finit-priority" }
            description       "This option controls the global compiler flags
                            which are used to compile all packages by default.
                            Individual packages may define options which
                            override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-m5206e -g -nostdlib -Wl,--gc-sections -Wl,-static" }

            description       "This option controls the global linker flags.
                            Individual packages may define options which
                            override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "ROMRAM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define

            description       "This option enables the building of the GDB
                            stubs for the board. The common HAL controls
                            take care of most of the build process, but the
                            final conversion from ELF image to binary data is
                            handled by the platform CDL, allowing relocation
                            of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.srec : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -S -O srec $< $@
            }
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { (CYG_HAL_STARTUP == "RAM") ? "coldfire_m5272c3_ram" : \
                     (CYG_HAL_STARTUP == "ROMRAM") ? "coldfire_m5272c3_romram" : \
                                            "coldfire_m5272c3_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { (CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_coldfire_m5272c3_ram.ldi>" : \
                         (CYG_HAL_STARTUP == "ROMRAM") ? "<pkgconf/mlt_coldfire_m5272c3_romram.ldi>" : \
                                                    "<pkgconf/mlt_coldfire_m5272c3_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { (CYG_HAL_STARTUP == "RAM") ? "<pkgconf/mlt_coldfire_m5272c3_ram.h>" : \
                         (CYG_HAL_STARTUP == "ROMRAM") ? "<pkgconf/mlt_coldfire_m5272c3_romram.h>" : \
                                                    "<pkgconf/mlt_coldfire_m5272c3_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "GDB_stubs" }
        default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
        requires      { CYG_HAL_STARTUP == "RAM" }
        parent        CYGPKG_HAL_ROM_MONITOR

        description       "Support can be enabled for boot ROMs or ROM
                        monitors which contain GDB stubs. This support
                        changes various eCos semantics such as the encoding of
                        diagnostic output, and the overriding of hardware
                        interrupt vectors."
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "ROMRAM" }

        description       "Enable this option if this program is to be used as
                        a ROM monitor, i.e. applications will be loaded into
                        RAM on the board, and this ROM monitor may process
                        exceptions or interrupts generated from the
                        application. This enables features such as utilizing
                        a separate interrupt stack when exceptions are
                        generated."
    }
}
