# ====================================================================
#
#      hal_arm_mac7100.cdl
#
#      Freescale MAC7100 HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Nick Garnett <nickg@calivar.com>
## Copyright (C) 2006 eCosCentric Ltd
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Ilija Koco <ilijak@siva.com.mk>
# Contributors:   
# Date:           2006-02-03
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_MAC7100 {
    display       "Freescale MAC7100 variant HAL"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_mac7100.h
    include_dir   cyg/hal
    hardware
    description   "
        The MAC7100 HAL package provides the support needed to run
        eCos on Freescale MAC7100 based targets."

    compile       flash_security.S hal_diag.c mac7100_misc.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT
    implements    CYGINT_HAL_ARM_ARCH_ARM7
    implements    CYGINT_HAL_ARM_THUMB_ARCH
    implements    CYGINT_HAL_ARM_BIGENDIAN
    requires { CYGHWR_HAL_ARM_BIGENDIAN == 1 }

    # Let the architectural HAL see this variant's files
    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_IO_H"
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_ARCH_H"
    }

    cdl_option CYGHWR_HAL_ARM_MAC7100 {
        display        "MAC7100 variant used"
        flavor         data
        default_value  {"MAC7111"}
        legal_values   {"MAC7111" "MAC7121" "MAC7116" }
        description    "
            The MAC7100 microcontroller family has several variants,
            the main differences being the amount of on-chip SRAM,
            peripherals and their layout. This option allows the
            platform HALs to select the specific microcontroller being
            used."
    }

    cdl_option CYGHWR_HAL_ARM_MAC7100_FIQ {
        display       "handle FIQ as an IRQ"
        flavor        bool
        default_value 0
        description   "
            Enable this option if you need to handle FIQ interrupts in the
            normal way, i.e. a FIQ interrupt will be treated as a normal IRQ 
            using the highest priority
            "
    }

    cdl_option CYGHWR_HAL_ARM_MAC7100_INTC_FIQDEF {
        display       "Set FIQDEF"
        flavor        data
        default_value CYGHWR_HAL_ARM_MAC7100_FIQ ? 14 : 16
        legal_values 0 to 32
        description   "
            Set maximum level that shall be routed to IRQ.
            "
    }

    cdl_option CYGHWR_HAL_ARM_MAC7100_INTC_EMASK {
        display       "enable INTC to automatically handle CLMASK"
        flavor        data
        default_value 0x20
        legal_values 0x00 0x20
        description   "
            Enable this option if you need INTC to automatically mask 
            lower level IRQ.
            
            - 0x00 - disable
            - 0x20 - enable
            
            "
    }
}
