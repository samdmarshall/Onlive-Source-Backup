# ====================================================================
#
#      flash_at91.cdl
#
#      FLASH programming for devices with the Embedded Flash Controller 
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2006 eCosCentric LTD
## Copyright (C) 2006 Andrew Lunn <andrew.lunn@ascom.ch>
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      dmoseley
# Original data:  gthomas
# Contributors:   Andrew Lunn, Oliver Munz
# Date:           2000-10-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_AT91 {
    display       "at91 FLASH memory support"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH

    implements    CYGHWR_IO_FLASH_DEVICE

    include_dir   .
    description   "FLASH memory device support for at91 EFC"
    compile       at91_flash.c
    
    cdl_option    CYGBLD_DEV_FLASH_AT91_LOCKING {
        display       "Support block locking"
        default_value 1
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        description   "
            The driver will implement flash block locking when this
            option is enabled. Note that the device implements sector
            locking, not block locking, where sectors are bigger than
            blocks. So the sector which contains the block will be
            locked/unlocked

            WARNING: The errata says that these lock bits only have 
            a life of 100 cycles for the AT91SAM7S devices."
    }
}

