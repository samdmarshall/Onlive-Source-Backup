# ====================================================================
#
#      ezxml.cdl
#
#      XML parser
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2005 eCosCentric Ltd
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Matt Jerdonek
# Original data:  Matt Jerdonek
# Contributors:
# Date:           2005-01-31
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_EZXML {
        display      "ezXML XML parser"
        description  "
            ezXML is a C library for parsing XML documents inspired by
            simpleXML for PHP.  As the name implies, it's easy to
            use. It's ideal for parsing xml configuration files or
            REST web service responses. It's also fast and lightweight
            (11k compiled)."

        compile      ezxml.c

        cdl_option CYGPKG_EZXML_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D__ECOS__" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are used in addition
                to the set of global flags."
        }
        
        cdl_option CYGPKG_EZXML_TESTS {
            display "ezXML tests"
            flavor  data
            no_define
            calculated { "tests/ezxml" }
        }
}
